entity cla is port(
    a, b : in std_logic_vector(7 downto 0);
    cin : in std_logic;
    s : out std_logic_vector(7 downto 0);
    cout : out std_logic;
);

architecture structural of cla is

    begin

        

end structural;