library ieee;
use ieee.std_logic_1164.all;

entity rotateleft is
    port(   
    	    a: in   std_logic_vector (7 downto 0);
    	    b: out  std_logic_vector (7 downto 0)
   	);
end rotateleft;
